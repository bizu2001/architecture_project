//this code , as a whole , follows the structure of the 65th page of PPT5. I have added pipeline to the design
//Please check the mentioned page if you could not understand my code
`timescale 100fs/100fs

//the pc register
module PC(clk,enable,next_pc,pc);
input clk;
input enable;
input[31:0] next_pc;
output reg[31:0] pc;
initial
begin
	pc=32'b00000000000000000000000000000000;
end
always@(posedge clk)
begin
	if(enable)
	begin
		pc<=next_pc;
	end

end
endmodule

//the instruction memory
module InstructionRAM
    ( // Inputs
      input  CLOCK // clock
    , input  ENABLE
    , input [31:0] FETCH_ADDRESS

      // Outputs
    , output  reg [31:0] DATA

    );
  // blockRamFile begin
  reg [31:0] RAM [0:512-1];

  initial begin
    $readmemb("instructions.bin",RAM);

  end
//  assign address = FETCH_ADDRESS/4;
always@(*) begin
if(ENABLE==1)
begin
 DATA = RAM[FETCH_ADDRESS/4];
end
end
endmodule
module MainMemory
    ( // Inputs
      input  CLOCK // clock
    , input  ENABLE
    , input [31:0] FETCH_ADDRESS
	, input [31:0] MEM_instruction
	, input memread
	, input memwrite
	, input [31:0]writedata

      // Outputs
    , output reg [31:0] DATA
    );
 

  // blockRam begin
  reg [31:0] DATA_RAM [0:512-1];

  reg [16383:0] ram_init;
  integer i;
  initial begin
    ram_init = {32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000,32'b00000000000000000000000000000000};
    for (i=0; i < 512; i = i + 1) begin
      DATA_RAM[512-1-i] = ram_init[i*32+:32];
    end
  end
 
  integer out_file;
  initial
  begin
	  out_file=$fopen("output.txt","w");
  end
  always@(*)begin
	  if(memwrite&ENABLE)
 	  begin
 		  DATA_RAM[FETCH_ADDRESS] =writedata;
 	  end
 	  if (memread&ENABLE)
 	  begin
 		  DATA = DATA_RAM[FETCH_ADDRESS];
 	  end
	  if(MEM_instruction == 32'b11111111111111111111111111111111)
	  begin
	  for(i=0;i<512;i=i+1)
	  begin
		  $display("the memory result is now stored in output.txt");
		  $display(DATA_RAM[i]);
		  $fwrite(out_file,"%b\n",DATA_RAM[i]);
	  end
	  end
  end
endmodule
//the IF/ID register
module IFIDreg(clk,en,IF_instruction,IF_pc,ID_pc,ID_instruction);
input clk,en;
input [31:0]IF_instruction;
input [31:0] IF_pc;
output reg[31:0] ID_pc;
output reg[31:0] ID_instruction;
always@(posedge clk)
begin
	if (en)
	begin
		ID_pc<=IF_pc;
		ID_instruction<=IF_instruction;
	end
end
endmodule
//the register file
//regwrite: enable to write in the register file
//a 32*32 register file
module registerfile(clk,readregister1,readregister2,writeregister,writedata,regwrite,readdata1,readdata2);
input clk;
input [4:0]readregister1;
input [4:0]readregister2;
input [4:0]writeregister;
input [31:0]writedata;
input regwrite;
output reg [31:0]readdata1;
output reg [31:0]readdata2;
reg[31:0] registers[31:0];
integer i;
initial
begin
	for(i=0;i<32;i++)
	begin
	registers[32-1-i]=32'b00000000000000000000000000000000;
	end
end
always@(posedge clk)
begin
	readdata1<=registers[readregister1];
	readdata2<=registers[readregister2];
	if(regwrite==1'b1)
	begin
		registers[writeregister]<=writedata;
	end
end
endmodule
//the control
//the control is a little different from that of PPT
//to simplify the process, alu control and control is combined!
module maincontrol(
input [5:0]opcode,
input [5:0]funct,
output reg[1:0] regdst,//add one bit to support jal operation(connect to the writeregsiter of the register file)
//regdet:01 from[15:11],00from [20:16],10from 11111
output reg regwrite,
output reg alusrc,
output reg [3:0] aluctr,
output reg pcsrc,
output reg memread,
output reg memwrite,
output reg [1:0]memtoreg,//add one bit to support jal,store pc+4 in the reg
//memtoreg:00from alu,01from mem, 10frompc+4
output reg jump,
output reg immctr,//whether zero extend or signextend for the imm
output reg jumpreg,//for jr
output reg pcbne);//determine the instruction is bne or beq
    always@(*)
    begin
        case(opcode)
        6'b000000:
        begin
            regdst<=2'b01;
			regwrite<=1'b1;
			alusrc<=1'b0;
            memread<=1'b0;
			memwrite<=1'b0;
			pcbne<=1'b0;
			pcsrc<=1'b0;
			immctr<=1'b0;
			jump<=1'b0;
			if (funct==001000)//jr
			begin
				aluctr<=4'b0000;
				memtoreg<=2'b00;
				jumpreg<=1'b1;
			end
			else
			begin
            memtoreg<=2'b00;
			jumpreg<=1'b0;
            case(funct)
                6'b100000://add
                begin
                    aluctr<=4'b0010;	
                end
                6'b100001://addu
                begin
                    aluctr<=4'b1011;
                end
                6'b100100://and
                begin
                    aluctr<=4'b0000;
                end
                6'b100010://sub
                begin
                    aluctr<=4'b0110;
                end
                6'b100011://subu
                begin
                    aluctr<=4'b1100;
                end
                6'b100101://or
                begin
                    aluctr<=4'b0001;
                end
                6'b100111://nor
                begin
                    aluctr<=4'b0011;
                end
                6'b100110://xor
                begin
                    aluctr<=4'b0100;
                end
                6'b000000://sll
                begin
                    aluctr<=4'b0101;
                end
                6'b000100://sllv
                begin
                    aluctr<=4'b1101;
                end
                6'b000010://srl
                begin
                    aluctr<=4'b0111;
                end
                6'b000110://srlv
                begin
                    aluctr<=4'b1110;
                end
                6'b000011://sra
                begin
                    aluctr<=4'b1000;
                end
                6'b000111://srav
                begin
                    aluctr<=4'b1111;
                end
                6'b101010://slt
                begin
                    aluctr<=4'b1001;
                end
                6'b101011://sltu
                begin
                    aluctr<=4'b1010;
                end
            endcase
		    end
        end
        6'b001010://slti
        begin
			regdst<=2'b00;
			regwrite<=1'b1;
            alusrc<=1'b1;
            aluctr<=4'b1001;//same as slt
            pcsrc<=1'b0;
			pcbne<=1'b0;
			memread<=1'b0;
			memwrite<=1'b0;
			memtoreg<=2'b00;
			jump<=1'b0;
			immctr<=1'b0;
			jumpreg<=1'b0;
        end
        6'b001011://sltiu
        begin
            alusrc<=1'b1;
            aluctr<=4'b1010;//same as sltu
			regdst<=2'b00;
			regwrite<=1'b1;
            pcsrc<=1'b0;
			pcbne<=1'b0;
			memread<=1'b0;
			memwrite<=1'b0;
			memtoreg<=2'b00;
			jump<=1'b0;
			immctr<=1'b0;
			jumpreg<=1'b0;
        end
        6'b100011://lw
        begin
            alusrc<=1'b1;
            aluctr<=4'b0010;//same as add
			regdst<=2'b00;
			regwrite<=1'b1;
            pcsrc<=1'b0;
			pcbne<=1'b0;
			memread<=1'b1;//load
			memwrite<=1'b0;
			memtoreg<=2'b01;//load
			jump<=1'b0;
			immctr<=1'b0;
			jumpreg<=1'b0;
        end
        6'b101011://sw
        begin
            alusrc<=1'b1;
            aluctr<=4'b0010;//same as add
			regdst<=2'b00;
			regwrite<=1'b0;//no need to write register
            pcsrc<=1'b0;
			pcbne<=1'b0;
			memread<=1'b0;
			memwrite<=1'b1;//save
			memtoreg<=2'b00;//don't care
			jump<=1'b0;
			immctr<=1'b0;
			jumpreg<=1'b0;
        end
        6'b000100://beq
        begin
            alusrc<=1'b0;
            aluctr<=4'b0110;//same as sub
			regdst<=2'b00;//don't care
			regwrite<=1'b0;
            pcsrc<=1'b1;//branch
			pcbne<=1'b1;//beq
			memread<=1'b0;//
			memwrite<=1'b0;
			memtoreg<=2'b00;//don't care
			jump<=1'b0;
			immctr<=1'b0;
			jumpreg<=1'b0;
        end
        6'b000101://bne
        begin
            alusrc<=1'b0;
            aluctr<=4'b0110;//same as sub
			regdst<=2'b00;//don't care
			regwrite<=1'b0;
            pcsrc<=1'b1;//branch
			pcbne<=1'b0;//bne
			memread<=1'b0;//
			memwrite<=1'b0;
			memtoreg<=2'b00;//don't care
			jump<=1'b0;
			immctr<=1'b0;
			jumpreg<=1'b0;
        end
        6'b001101://ori
        begin
            alusrc<=1'b1;
            aluctr<=4'b0001;
			regdst<=2'b00;
			regwrite<=1'b1;
            pcsrc<=1'b0;
			pcbne<=1'b0;
			memread<=1'b0;
			memwrite<=1'b0;
			memtoreg<=2'b00;
			jump<=1'b0;
			immctr<=1'b1;//zero extend
			jumpreg<=1'b0;
        end
        6'b001100://andi
        begin
            alusrc<=1'b1;
            aluctr<=4'b0000;
			regdst<=2'b00;
			regwrite<=1'b1;
            pcsrc<=1'b0;
			pcbne<=1'b0;
			memread<=1'b0;
			memwrite<=1'b0;
			memtoreg<=2'b00;
			jump<=1'b0;
			immctr<=1'b1;//zero extend
			jumpreg<=1'b0;
        end
        6'b001110://xori
        begin
            alusrc<=1'b1;
            aluctr<=4'b0100;
			regdst<=2'b00;
			regwrite<=1'b1;
            pcsrc<=1'b0;
			pcbne<=1'b0;
			memread<=1'b0;
			memwrite<=1'b0;
			memtoreg<=2'b00;
			jump<=1'b0;
			immctr<=1'b1;//zero extend
			jumpreg<=1'b0;
        end
        6'b001000://addi
        begin
            alusrc<=1'b1;
            aluctr<=4'b0010;//same as add
			regdst<=2'b00;
			regwrite<=1'b1;
            pcsrc<=1'b0;
			pcbne<=1'b0;
			memread<=1'b0;
			memwrite<=1'b0;
			memtoreg<=2'b00;
			jump<=1'b0;
			immctr<=1'b0;//sign extend
			jumpreg<=1'b0;
        end
        6'b001001://addiu
        begin
            alusrc<=1'b1;
            aluctr<=4'b1011;//same as addu
			regdst<=2'b00;
			regwrite<=1'b1;
            pcsrc<=1'b0;
			pcbne<=1'b0;
			memread<=1'b0;
			memwrite<=1'b0;
			memtoreg<=2'b00;
			jump<=1'b0;
			immctr<=1'b0;//sign extend
			jumpreg<=1'b0;
        end
		6'b000010://j
		begin
			alusrc<=1'b1;//don't care
            aluctr<=4'b0000;//don't care
			regdst<=2'b00;//don't care
			regwrite<=1'b0;
            pcsrc<=1'b0;//don't care
			pcbne<=1'b0;//don't care
			memread<=1'b0;
			memwrite<=1'b0;
			memtoreg<=2'b00;//don't care
			jump<=1'b1;
			immctr<=1'b0;//don't care
			jumpreg<=1'b0;
		end
		6'b000011://jal
		begin
			alusrc<=1'b1;//don't care
            aluctr<=4'b0000;//don't care
			regdst<=2'b10;//number 11111
			regwrite<=1'b1;
            pcsrc<=1'b0;//don't care
			pcbne<=1'b0;//don't care
			memread<=1'b0;
			memwrite<=1'b0;
			memtoreg<=2'b10;//return pc+4
			jump<=1'b1;
			immctr<=1'b0;//don't care
			jumpreg<=1'b0;
		end
		default:
		begin
			alusrc<=1'b0;
            aluctr<=4'b0000;
			regdst<=2'b00;
			regwrite<=1'b0;
            pcsrc<=1'b0;
			pcbne<=1'b0;
			memread<=1'b0;
			memwrite<=1'b0;
			memtoreg<=2'b00;
			jump<=1'b0;
			immctr<=1'b0;
			jumpreg<=1'b0;
		end	
        endcase
    end
endmodule

module imm(imm,immctr,immoper);//sign extend the 16 bits imm
input [15:0]imm;
input immctr;
output reg[31:0] immoper;
always@(*)
begin
	if (immctr==1'b0)
	begin
		immoper = {{16{imm[15]}},imm};
	end
	if (immctr==1'b1)
	begin
		immoper = {{16{1'b0}},imm};
	end
end
endmodule

module IDEXreg(input clk, input en,input [31:0]IDreaddata1,input[31:0]IDreaddata2,
input [31:0]IDimmoper,input [1:0]IDregdst,input [3:0]IDaluctr,input IDalusrc,input IDregwrite,
input IDpcsrc,input IDpcbne,input IDmemread,input IDmemwrite,input [1:0]IDmemtoreg,
input IDjump,input IDjumpreg,input [31:0]IDPC,input [31:0] shamt,input [4:0]IDins2016,input [4:0]IDins1511,
input [25:0]IDjumpimm,input [31:0]ID_instruction,output reg[31:0] EXreaddata1,output reg[31:0] EXreaddata2,output reg[31:0] EXimmoper,
output reg[3:0]EXaluctr,output reg EXalusrc,output reg[1:0]EXregdst,
output reg EXregwrite,output reg EXpcsrc,output reg EXpcbne,
output reg EXmemread,output reg EXmemwrite,output reg[1:0]EXmemtoreg,
output reg EXjump,output reg EXjumpreg, output reg[31:0]EXPC, output reg[31:0] EXshamt,
output reg[4:0] EXins2016,output reg[4:0] EXins1511,output reg[25:0]EXjumpimm, output reg[31:0]EX_instruction);
always@(posedge clk)
begin
	if (en)
	begin
		EXreaddata1<=IDreaddata1;
		EXreaddata2<=IDreaddata2;
		EXimmoper<=IDimmoper;
		EXaluctr<=IDaluctr;
		EXalusrc<=IDalusrc;
		EXregdst<=IDregdst;
		EXregwrite<=IDregwrite;
		EXpcsrc<=IDpcsrc;
		EXpcbne<=IDpcbne;
		EXmemread<=IDmemread;
		EXmemwrite<=IDmemwrite;
		EXmemtoreg<=IDmemtoreg;
		EXjump<=IDjump;
		EXjumpreg<=IDjumpreg;
		EXPC<=IDPC;
		EXshamt<=shamt;
		EXins2016<=IDins2016;
		EXins1511<=IDins1511;
		EXjumpimm<=IDjumpimm;
		EX_instruction<=ID_instruction;
	end
end
endmodule

module ALU(aluctr,A,B,shamt,result,zero,overflow);
input[31:0] A;
input[31:0] B;
input [3:0] aluctr;
input [31:0] shamt;
output reg[31:0] result;
output  reg zero;
output  reg overflow;
always@(*)begin
    case(aluctr)
    4'b0010://add
    begin
        result = A+B;
        overflow = (A[31]^B[31]) ? 0: (result[31]^A[31]);
        zero = result?0:1;
    end
    4'b1011://addu
    begin
        result = A+B;
        overflow =1'b0;
        zero = result?0:1;
    end
    4'b0000://and
    begin
        result = A&B;
        overflow =1'b0;
        zero = result?0:1;
    end
    4'b0110://sub
    begin
        result = $signed(A)-$signed(B);
        overflow = (A[31]^B[31]) ? (result[31]^A[31]):0;
        zero = result?0:1;
    end
    4'b1100://subu
    begin
        result=$signed(A)-$signed(B);
        overflow =1'b0;
        zero = result?0:1;
    end
    4'b0001://or
    begin
        result = A|B;
        overflow =1'b0;
        zero = result?0:1;
    end
    4'b0011://nor
    begin
        result=~(A|B);
        overflow =1'b0;
        zero = result?0:1;
    end
    4'b0100://xor
    begin
        result = A^B;
        overflow =1'b0;
        zero = result?0:1;
    end
    4'b0101://sll
    begin
        result=B<<shamt[4:0];
        overflow =1'b0;
        zero = result?0:1;
    end
    4'b1101://sllv
    begin
        result=B<<A[4:0];
        overflow =1'b0;
        zero = result?0:1;
    end
    4'b0111://srl
    begin
        result=B>>shamt[4:0];
        overflow =1'b0;
        zero = result?0:1;
    end
    4'b1110://srlv
    begin
        result=B>>A[4:0];
        overflow =1'b0;
        zero = result?0:1;
    end
    4'b1000://sra
    begin
        result = $signed($signed(B) >>> shamt[4:0]);
        overflow =1'b0;
        zero = result?0:1;
    end
    4'b1111://srav
    begin
        result = $signed($signed(B) >>> A[4:0]);
        overflow =1'b0;
        zero = result?0:1;
    end
    4'b1001://slt
    begin
        result=($signed(A)<$signed(B))?32'b1:32'b0;
        overflow =1'b0;
        zero = result?0:1;
    end
    4'b1010://sltu
    begin
        result = (A<B) ? 32'b1 : 32'b0;
        overflow =1'b0;
        zero = result?0:1;
    end
    endcase
end
endmodule

//adder will return the value of a and b
module adder(a,b,result);
input [31:0]a;
input [31:0]b;
output reg[31:0]result;
always@(*)
begin
	result=a+b;
end
endmodule

//the EX/MEM pipeline
module EXMEMreg(input clk, input en,
input EXregwrite,input EXpcsrc,input EXpcbne,input EXmemread,
input EXmemwrite,input [1:0]EXmemtoreg,input EXjump,input EXjumpreg, input [31:0]EXPC_A,//EXPC_A = EXPC
input [31:0]EXIPC,input EXzero, input [31:0]EXresult,input [31:0]EXreaddata1,//EXIPC=EXPC+immoper<<2
input [31:0]EXreaddata2,input [4:0]EXdst,input [31:0]EXjumpadd, input [31:0] EX_instruction, output reg MEMregwrite, output reg MEMpcsrc,
output reg MEMpcbne, output reg MEMmemread, output reg MEMmemwrite, output reg[1:0]MEMmemtoreg,
output reg MEMjump,output reg MEMjumpreg,output reg [31:0]MEMPC_A,output reg[31:0]MEMPC, output reg MEMzero,
output reg[31:0] MEMresult,output reg [31:0]MEMreaddata1,
output reg [31:0]MEMreaddata2, output reg[4:0]MEMdst,output reg[31:0]MEMjumpadd,output reg[31:0]MEM_instruction);
always@(posedge clk)
begin
	if (en)
	begin
		MEMregwrite<=EXregwrite;
		MEMpcsrc<=EXpcsrc;
        MEMpcbne<=EXpcbne;
		MEMmemread<=EXmemread;
		MEMmemwrite<=EXmemwrite;
		MEMmemtoreg<=EXmemtoreg;
		MEMjump<=EXjump;
		MEMjumpreg<=EXjumpreg;
		MEMPC_A<=EXPC_A;
		MEMPC<=EXIPC;
		MEMzero<=EXzero;
		MEMresult<=EXresult;
		MEMreaddata1<=EXreaddata1;
		MEMreaddata2<=EXreaddata2;
		MEMdst<=EXdst;
		MEMjumpadd<=EXjumpadd;
		MEM_instruction<=EX_instruction;
	end
		
end
endmodule

module MEMWBreg(input clk, input en, input MEMregwrite,input [1:0]MEMmemtoreg,
input [31:0]MEMreaddata, input [31:0]MEMresult, input [4:0]MEMdst,input [31:0]MEMPC_A,output reg WBregwrite,
output reg[1:0] WBmemtoreg, output reg[31:0] WBreaddata, output reg[31:0]WBresult,
output reg[4:0] WBdst,output reg[31:0]WBPC);
always@(posedge clk)
begin
	if(en)
	begin
		WBregwrite<=MEMregwrite;
		WBmemtoreg<=MEMmemtoreg;
		WBreaddata<=MEMreaddata;
		WBresult<=MEMresult;
		WBdst<=MEMdst;
	end
end
endmodule

// module hazardunit();

// endmodule

module twoMUX(a,b,sel,out);//if sel = 0,choose a;
input [31:0] a;
input [31:0] b;
input sel;
output reg[31:0]out;
always@(*)
begin
out = sel?b:a;
end
endmodule

module threeMUX32(a,b,c,sel,out);//a:00,b:01,c:10
input [31:0] a;
input [31:0] b;
input [31:0] c;
input [1:0]sel;
output reg[31:0]out;
always@(*)
begin
out = sel[1] ? c: (sel[0]? b : a); 
end
endmodule

module threeMUX5(a,b,c,sel,out);//a:00,b:01,c:10
input [4:0] a;
input [4:0] b;
input [4:0] c;
input [1:0]sel;
output reg[4:0]out;
always@(*)
begin
 out = sel[1] ? c: (sel[0]? b : a); 
end
endmodule

module CPU(clk);
input clk;
// clk clock(enable,clk);
wire [31:0] pc;
wire enable = 1'b1;
wire [31:0] IF_pc;
wire [31:0] IF_instruction;
wire [31:0] ID_pc;
wire [31:0] ID_instruction;

PC programcounter(clk,enable,next_pc,pc);
adder adder1(pc,32'b00000000000000000000000000000100,IF_pc);//IF_pc = pc+4;
InstructionRAM instructionfile(clk,enable,pc,IF_instruction);
IFIDreg pipeline1(clk,enable,IF_instruction,IF_pc,ID_pc,ID_instruction);
//the ID stage
wire [5:0] opcode;
wire [5:0] funct;
wire [4:0] rs;
wire [4:0] rt;
wire [15:0] imm;
wire [31:0] shamt;
wire [4:0] IDins2016;
wire [4:0] IDins1511;
wire [25:0] IDjumpimm;

assign opcode = ID_instruction[31:26];
assign funct = ID_instruction[5:0];
assign rs = ID_instruction[25:21];
assign rt = ID_instruction[20:16];
assign imm = ID_instruction[15:0];
assign shamt = {{27{1'b0}},ID_instruction[10:6]};
assign IDins2016 = ID_instruction[20:16];
assign IDins1511 = ID_instruction[15:11];
assign IDjumpimm = ID_instruction[25:0];

wire [1:0] regdst;
wire regwrite;
wire alusrc;
wire [3:0] aluctr;
wire pcsrc;
wire memread;
wire memwrite;
wire [1:0] memtoreg;
wire jump;
wire immctr;
wire jumpreg;
wire pcbne;
wire [31:0] IDimmoper;
maincontrol control(opcode,funct,regdst,
regwrite,alusrc,aluctr,pcsrc,memread,memwrite,memtoreg,jump,
immctr,jumpreg,pcbne);
imm immextender(imm,immctr,IDimmoper);//IDimmoper is the sign extended imm 
wire [31:0] IDreaddata1;
wire [31:0] IDreaddata2;
registerfile regfile(clk,rs,rt,WBdst,WBwritedata,WBregwrite,IDreaddata1,IDreaddata2);
wire [31:0] EXreaddata1;
wire [31:0] EXreaddata2;
wire [31:0] EXimmoper;
wire [3:0] EXaluctr;
wire EXalusrc;
wire [1:0] EXregdst;
wire EXregwrite;
wire EXpcsrc;
wire EXpcbne;
wire EXmemread;
wire EXmemwrite;
wire [1:0]EXmemtoreg;
wire EXjump;
wire EXjumpreg;
wire [31:0]EXPC;
wire [31:0]EXshamt;
wire [4:0] EXins2016;
wire [4:0] EXins1511;
wire [25:0] EXjumpimm;
wire [31:0] EX_instruction;
IDEXreg pipeline2(clk,enable,IDreaddata1,IDreaddata2,
IDimmoper,regdst,aluctr,alusrc,regwrite,
pcsrc,pcbne,memread,memwrite,memtoreg,
jump,jumpreg,ID_pc,shamt,IDins2016,IDins1511,IDjumpimm,ID_instruction,
EXreaddata1,EXreaddata2,EXimmoper,
EXaluctr,EXalusrc,EXregdst,
EXregwrite,EXpcsrc,EXpcbne,
EXmemread,EXmemwrite,EXmemtoreg,
EXjump, EXjumpreg, EXPC,EXshamt,
EXins2016,EXins1511,EXjumpimm,EX_instruction);
//EX stage
wire [31:0] EXIPC;
adder adder2(EXPC,EXimmoper<<2,EXIPC);
wire [31:0]EXjumpadd;
assign EXjumpadd = {{EXPC[31:28]},{EXjumpimm},{2'b00}};//the jump address
wire [31:0]B;
twoMUX mux1(EXreaddata2,EXimmoper,EXalusrc,B);//B is the second input to the ALU
wire [31:0] result;
wire zero;
wire overflow;
ALU ALU(EXaluctr,EXreaddata1,B,EXshamt,result,zero,overflow);//EXreaddata1 is the first input to the ALU, 
wire [4:0] EXdst;
threeMUX5 mux2(EXins2016,EXins1511,5'b11111,EXregdst,EXdst);
wire MEMregwrite;
wire MEMpcsrc;
wire MEMpcbne;
wire MEMmemread;
wire MEMmemwrite;
wire [1:0] MEMmemtoreg;
wire MEMjump;
wire MEMjumpreg;
wire [31:0]MEMPC_A;
wire [31:0]MEMPC;
wire MEMzero;
wire [31:0] MEMresult;
wire [31:0] MEMreaddata1;
wire [31:0] MEMreaddata2;
wire [4:0] MEMdst;
wire [31:0] MEMjumpadd;
wire [31:0] MEM_instruction;
EXMEMreg pipeline3(clk, enable,EXregwrite,EXpcsrc,EXpcbne,
EXmemread,EXmemwrite,EXmemtoreg,EXjump,
EXjumpreg,EXPC ,EXIPC,zero, result,EXreaddata1,
EXreaddata2,EXdst,EXjumpadd,EX_instruction, MEMregwrite, MEMpcsrc,
MEMpcbne, MEMmemread,MEMmemwrite, MEMmemtoreg,
MEMjump,MEMjumpreg,MEMPC_A,MEMPC, MEMzero,
MEMresult,MEMreaddata1,MEMreaddata2, MEMdst,MEMjumpadd,MEM_instruction);
wire [31:0]MEMReadData;
MainMemory MainMemory(clk,enable,MEMresult,MEM_instruction, MEMmemread,
MEMmemwrite,MEMreaddata2,MEMReadData);
wire branch;
wire [31:0]out1;
wire [31:0]out2;
wire [31:0]next_pc;
assign branch = MEMpcsrc&(~pcbne^MEMzero);
twoMUX mux3(IF_pc,MEMPC,branch,out1);//select the next pc: branch address or pc+4
twoMUX mux4(out1,MEMjumpadd,MEMjump,out2);//select the next pc: whether to use jump address
twoMUX mux5(out2,MEMreaddata1,MEMjumpreg,next_pc);//select the next pc: whether to jump to the address in the regsiter(jr)
//WB stage
wire WBregwrite;
wire [1:0]WBmemtoreg;
wire [31:0]WBreaddata;
wire [31:0]WBresult;
wire  [4:0]WBdst;
wire [31:0]WBPC;
MEMWBreg pipeline4(clk, enable,MEMregwrite,MEMmemtoreg,
MEMReadData, MEMresult, MEMdst,MEMPC_A,WBregwrite,
WBmemtoreg, WBreaddata, WBresult,
WBdst,WBPC);
wire[31:0]WBwritedata;//WBdata is the data that will write back to the register file
threeMUX32 mux6(WBresult,WBreaddata,WBPC,WBmemtoreg,WBwritedata);

endmodule


 